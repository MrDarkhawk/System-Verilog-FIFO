////////////////////////////////////////////////
//
//           HEADER
//
/////////////////////////////////////////////////

`ifndef FIFO_DEFINES_SV
`define FIFO_DEFINES_SV

`define ADDR_WIDTH 4
`define DATA_WIDTH 8

`endif